----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:56:41 05/18/2022 
-- Design Name: 
-- Module Name:    PromedioB - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PromedioB is
	Port(A, B : IN STD_LOGIC_VECTOR (0 TO 3);
			C: OUT STD_LOGIC_VECTOR (0 TO 3));
end PromedioB;

architecture Behavioral of PromedioB is

begin


end Behavioral;

