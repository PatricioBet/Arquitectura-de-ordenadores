----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:41:02 05/18/2022 
-- Design Name: 
-- Module Name:    circuitoFlujoDatosVector - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity circuitoFlujoDatosVector is
           port(a, b : in  STD_LOGIC_VECTOR (0 TO 3);
           F : in  STD_LOGIC);
end circuitoFlujoDatosVector;

architecture Behavioral of circuitoFlujoDatosVector is

begin


end Behavioral;

