----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:46:15 05/18/2022 
-- Design Name: 
-- Module Name:    promedioA - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity promedioA is
	Port(A, B : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			C: OUT STD_LOGIC_VECTOR (2 DOWNTO 0));
end PromedioA;

architecture Behavioral of promedioA is

begin


end Behavioral;

