----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:53:28 05/18/2022 
-- Design Name: 
-- Module Name:    Promedio - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

--ejercicio 1.11 a

entity Promedio is
Port(A, B : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			C: OUT STD_LOGIC_VECTOR (2 DOWNTO 0));
end Promedio;

architecture Behavioral of Promedio is

begin


end Behavioral;

